library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- initializing all sprites
-- sprite size: 16x16

entity Sprites is
   port(
      address	: in std_logic_vector(7 downto 0);
      dataOut	: out std_logic_vector(15 downto 0)
   );
end Sprites;

architecture Behavioral of Sprites is

type array_atom is array (15 downto 0) of std_logic_vector(15 downto 0); 
--constant ROM: array_atom:=(
signal symbol_player : array_atom; 
signal symbol_wall	: array_atom; 
signal symbol_0		: array_atom; --to display the scores/level
signal symbol_1		: array_atom;
signal symbol_2		: array_atom;
signal symbol_3		: array_atom; 
signal symbol_4		: array_atom;
signal symbol_5		: array_atom;
signal symbol_6		: array_atom; 
signal symbol_7		: array_atom;
signal symbol_8		: array_atom;
signal symbol_9		: array_atom; 
signal symbol_S		: array_atom; --todisplay the word scores
signal symbol_C		: array_atom;
signal symbol_O		: array_atom; 
signal symbol_R		: array_atom;
signal symbol_E		: array_atom;
signal symbol_L		: array_atom; -- to display the word LEVEL
signal symbol_V		: array_atom;

symbol_player( 0) <= "1111111111111111"; 
symbol_player( 1) <= "1100000000000011"; 
symbol_player( 2) <= "1100000000000011"; 
symbol_player( 3) <= "1101111001111011"; 
symbol_player( 4) <= "1100011001100011"; 
symbol_player( 5) <= "1100000000000011"; 
symbol_player( 6) <= "1100000000000011"; 
symbol_player( 7) <= "1100000000000011"; 
symbol_player( 8) <= "1100011111100011"; 
symbol_player( 9) <= "1100001111000011"; 
symbol_player(10) <= "1100000110000011"; 
symbol_player(11) <= "1100000000000011"; 
symbol_player(12) <= "1100000000000011"; 
symbol_player(13) <= "1100000000000011"; 
symbol_player(14) <= "1100000000000011";
symbol_player(15) <= "1100000000000011"; 
 
symbol_wall( 0) <= "1111111111111111"; 
symbol_wall( 1) <= "1001001001001001"; 
symbol_wall( 2) <= "1010010010010011"; 
symbol_wall( 3) <= "1100100100100101"; 
symbol_wall( 4) <= "1001001001001001"; 
symbol_wall( 5) <= "1010010010010011"; 
symbol_wall( 6) <= "1100100100100101"; 
symbol_wall( 7) <= "1001001001001001"; 
symbol_wall( 8) <= "1010010010010011"; 
symbol_wall( 9) <= "1100100100100101"; 
symbol_wall(10) <= "1001001001001001"; 
symbol_wall(11) <= "1010010010010011"; 
symbol_wall(12) <= "1100100100100101"; 
symbol_wall(13) <= "1001001001001001"; 
symbol_wall(14) <= "1010010010010011"; 
symbol_wall(15) <= "1111111111111111";  
 
symbol_L( 0) <= "0000000000000000";
symbol_L( 1) <= "0000000000000000";
symbol_L( 2) <= "0000000000000000";
symbol_L( 3) <= "0001100000000000";
symbol_L( 4) <= "0001100000000000";
symbol_L( 5) <= "0001100000000000";
symbol_L( 6) <= "0001100000000000";
symbol_L( 7) <= "0001100000000000";
symbol_L( 8) <= "0001100000000000";
symbol_L( 9) <= "0001100000000000";
symbol_L(10) <= "0001100000000000";
symbol_L(11) <= "0001111111111000";
symbol_L(12) <= "0001111111111000";
symbol_L(13) <= "0000000000000000";
symbol_L(14) <= "0000000000000000";
symbol_L(15) <= "0000000000000000";

symbol_V( 0) <= "0000000000000000";
symbol_V( 1) <= "0000000000000000";
symbol_V( 2) <= "0000000000000000";
symbol_V( 3) <= "0011000000001100";
symbol_V( 4) <= "0011000000001100";
symbol_V( 5) <= "0001100000011000";
symbol_V( 6) <= "0001100000011000";
symbol_V( 7) <= "0000110000110000";
symbol_V( 8) <= "0000110000011000";
symbol_V( 9) <= "0000011000110000";
symbol_V(10) <= "0000001111000000";
symbol_V(11) <= "0000000110000000";
symbol_V(12) <= "0000000000000000";
symbol_V(13) <= "0000000000000000";
symbol_V(14) <= "0000000000000000";
symbol_V(15) <= "0000000000000000";
 
symbol_S( 0) <= "0000000000000000";
symbol_S( 1) <= "0000000000000000";
symbol_S( 2) <= "0000000000000000";
symbol_S( 3) <= "0000111111111000";
symbol_S( 4) <= "0001111111111000";
symbol_S( 5) <= "0001100000000000";
symbol_S( 6) <= "0001100000000000";
symbol_S( 7) <= "0001111111111000";
symbol_S( 8) <= "0000111111111000";
symbol_S( 9) <= "0000000000011000";
symbol_S(10) <= "0000000000011000";
symbol_S(11) <= "0001111111111000";
symbol_S(12) <= "0001111111110000";
symbol_S(13) <= "0000000000000000";
symbol_S(14) <= "0000000000000000";
symbol_S(15) <= "0000000000000000";

symbol_C( 0) <= "0000000000000000";
symbol_C( 1) <= "0000000000000000";
symbol_C( 2) <= "0000000000000000";
symbol_C( 3) <= "0000111111111000";
symbol_C( 4) <= "0001111111111000";
symbol_C( 5) <= "0001100000000000";
symbol_C( 6) <= "0001100000000000";
symbol_C( 7) <= "0001100000000000";
symbol_C( 8) <= "0001100000000000";
symbol_C( 9) <= "0001100000000000";
symbol_C(10) <= "0001100000000000";
symbol_C(11) <= "0001111111111000";
symbol_C(12) <= "0000111111111000";
symbol_C(13) <= "0000000000000000";
symbol_C(14) <= "0000000000000000";
symbol_C(15) <= "0000000000000000";

symbol_O( 0) <= "0000000000000000";
symbol_O( 1) <= "0000000000000000";
symbol_O( 2) <= "0000000000000000";
symbol_O( 3) <= "0000111111110000";
symbol_O( 4) <= "0001111111111000";
symbol_O( 5) <= "0001100000011000";
symbol_O( 6) <= "0001100000011000";
symbol_O( 7) <= "0001100000011000";
symbol_O( 8) <= "0001100000011000";
symbol_O( 9) <= "0001100000011000";
symbol_O(10) <= "0001100000011000";
symbol_O(11) <= "0001111111111000";
symbol_O(12) <= "0000111111110000";
symbol_O(13) <= "0000000000000000";
symbol_O(14) <= "0000000000000000";
symbol_O(15) <= "0000000000000000";

symbol_R( 0) <= "0000000000000000";
symbol_R( 1) <= "0000000000000000";
symbol_R( 2) <= "0000000000000000";
symbol_R( 3) <= "0000111111110000";
symbol_R( 4) <= "0001111111111000";
symbol_R( 5) <= "0001100000011000";
symbol_R( 6) <= "0001100000011000";
symbol_R( 7) <= "0001111111111000";
symbol_R( 8) <= "0001111111110000";
symbol_R( 9) <= "0001100111000000";
symbol_R(10) <= "0001100011100000";
symbol_R(11) <= "0001100001110000";
symbol_R(12) <= "0001100000111000";
symbol_R(13) <= "0000000000000000";
symbol_R(14) <= "0000000000000000";
symbol_R(15) <= "0000000000000000";

symbol_E( 0) <= "0000000000000000";
symbol_E( 1) <= "0000000000000000";
symbol_E( 2) <= "0000000000000000";
symbol_E( 3) <= "0001111111111000";
symbol_E( 4) <= "0001111111111000";
symbol_E( 5) <= "0001100000000000";
symbol_E( 6) <= "0001100000000000";
symbol_E( 7) <= "0001111111111000";
symbol_E( 8) <= "0001111111111000";
symbol_E( 9) <= "0001100000000000";
symbol_E(10) <= "0001100000000000";
symbol_E(11) <= "0001111111111000";
symbol_E(12) <= "0001111111111000";
symbol_E(13) <= "0000000000000000";
symbol_E(14) <= "0000000000000000";
symbol_E(15) <= "0000000000000000";

symbol_0( 0) <= "0000000000000000";
symbol_0( 1) <= "0000000000000000";
symbol_0( 2) <= "0000000000000000";
symbol_0( 3) <= "0000111111110000";
symbol_0( 4) <= "0001111111111000";
symbol_0( 5) <= "0001100000011000";
symbol_0( 6) <= "0001100000011000";
symbol_0( 7) <= "0001100000011000";
symbol_0( 8) <= "0001100000011000";
symbol_0( 9) <= "0001100000011000";
symbol_0(10) <= "0001100000011000";
symbol_0(11) <= "0001111111111000";
symbol_0(12) <= "0000111111110000";
symbol_0(13) <= "0000000000000000";
symbol_0(14) <= "0000000000000000";
symbol_0(15) <= "0000000000000000";

symbol_1( 0) <= "0000000000000000";
symbol_1( 1) <= "0000000000000000";
symbol_1( 2) <= "0000000000000000";
symbol_1( 3) <= "0000001111000000";
symbol_1( 4) <= "0000011111000000";
symbol_1( 5) <= "0000111111000000";
symbol_1( 6) <= "0000000111000000";
symbol_1( 7) <= "0000000111000000";
symbol_1( 8) <= "0000000111000000";
symbol_1( 9) <= "0000000111000000";
symbol_1(10) <= "0000000111000000";
symbol_1(11) <= "0000000111000000";
symbol_1(12) <= "0000000111000000";
symbol_1(13) <= "0000000000000000";
symbol_1(14) <= "0000000000000000";
symbol_1(15) <= "0000000000000000";

symbol_2( 0) <= "0000000000000000";
symbol_2( 1) <= "0000000000000000";
symbol_2( 2) <= "0000000000000000";
symbol_2( 3) <= "0000111111110000";
symbol_2( 4) <= "0001111111111000";
symbol_2( 5) <= "0001110000111000";
symbol_2( 6) <= "0000000000111000";
symbol_2( 7) <= "0000000001110000";
symbol_2( 8) <= "0000000011100000";
symbol_2( 9) <= "0000000111000000";
symbol_2(10) <= "0000001110000000";
symbol_2(11) <= "0000111111111000";
symbol_2(12) <= "0001111111111000";
symbol_2(13) <= "0000000000000000";
symbol_2(14) <= "0000000000000000";
symbol_2(15) <= "0000000000000000";

symbol_3( 0) <= "0000000000000000";
symbol_3( 1) <= "0000000000000000";
symbol_3( 2) <= "0000000000000000";
symbol_3( 3) <= "0000111111110000";
symbol_3( 4) <= "0001111111111000";
symbol_3( 5) <= "0001100000011000";
symbol_3( 6) <= "0000000000011000";
symbol_3( 7) <= "0000000111110000";
symbol_3( 8) <= "0000000111110000";
symbol_3( 9) <= "0000000000011000";
symbol_3(10) <= "0001100000011000";
symbol_3(11) <= "0001111111111000";
symbol_3(12) <= "0000111111110000";
symbol_3(13) <= "0000000000000000";
symbol_3(14) <= "0000000000000000";
symbol_3(15) <= "0000000000000000";

symbol_4( 0) <= "0000000000000000";
symbol_4( 1) <= "0000000000000000";
symbol_4( 2) <= "0000000000000000";
symbol_4( 3) <= "0000000011111000";
symbol_4( 4) <= "0000000111111000";
symbol_4( 5) <= "0000001110011000";
symbol_4( 6) <= "0000011100011000";
symbol_4( 7) <= "0000111000011000";
symbol_4( 8) <= "0001111111111100";
symbol_4( 9) <= "0001111111111100";
symbol_4(10) <= "0000000000011000";
symbol_4(11) <= "0000000000011000";
symbol_4(12) <= "0000000000011000";
symbol_4(13) <= "0000000000000000";
symbol_4(14) <= "0000000000000000";
symbol_4(15) <= "0000000000000000";

symbol_5( 0) <= "0000000000000000";
symbol_5( 1) <= "0000000000000000";
symbol_5( 2) <= "0000000000000000";
symbol_5( 3) <= "0001111111111000";
symbol_5( 4) <= "0001111111111000";
symbol_5( 5) <= "0001100000000000";
symbol_5( 6) <= "0001100000000000";
symbol_5( 7) <= "0001111111110000";
symbol_5( 8) <= "0001111111111000";
symbol_5( 9) <= "0000000000011000";
symbol_5(10) <= "0001100000011000";
symbol_5(11) <= "0001111111111000";
symbol_5(12) <= "0000111111110000";
symbol_5(13) <= "0000000000000000";
symbol_5(14) <= "0000000000000000";
symbol_5(15) <= "0000000000000000";

symbol_6( 0) <= "0000000000000000";
symbol_6( 1) <= "0000000000000000";
symbol_6( 2) <= "0000000000000000";
symbol_6( 3) <= "0000111111110000";
symbol_6( 4) <= "0001111111111000";
symbol_6( 5) <= "0001100000011000";
symbol_6( 6) <= "0001100000000000";
symbol_6( 7) <= "0001111111110000";
symbol_6( 8) <= "0001111111111000";
symbol_6( 9) <= "0001100000011000";
symbol_6(10) <= "0001100000011000";
symbol_6(11) <= "0001111111111000";
symbol_6(12) <= "0000111111110000";
symbol_6(13) <= "0000000000000000";
symbol_6(14) <= "0000000000000000";
symbol_6(15) <= "0000000000000000";

symbol_7( 0) <= "0000000000000000";
symbol_7( 1) <= "0000000000000000";
symbol_7( 2) <= "0000000000000000";
symbol_7( 3) <= "0001111111111000";
symbol_7( 4) <= "0001111111111000";
symbol_7( 5) <= "0000000001110000";
symbol_7( 6) <= "0000000001110000";
symbol_7( 7) <= "0000000011100000";
symbol_7( 8) <= "0000000011100000";
symbol_7( 9) <= "0000000111000000";
symbol_7(10) <= "0000000111000000";
symbol_7(11) <= "0000001110000000";
symbol_7(12) <= "0000001110000000";
symbol_7(13) <= "0000000000000000";
symbol_7(14) <= "0000000000000000";
symbol_7(15) <= "0000000000000000";

symbol_8( 0) <= "0000000000000000";
symbol_8( 1) <= "0000000000000000";
symbol_8( 2) <= "0000000000000000";
symbol_8( 3) <= "0000111111110000";
symbol_8( 4) <= "0001111111111000";
symbol_8( 5) <= "0001100000011000";
symbol_8( 6) <= "0001100000011000";
symbol_8( 7) <= "0000111111110000";
symbol_8( 8) <= "0000111111110000";
symbol_8( 9) <= "0001100000011000";
symbol_8(10) <= "0001100000011000";
symbol_8(11) <= "0001111111111000";
symbol_8(12) <= "0000111111110000";
symbol_8(13) <= "0000000000000000";
symbol_8(14) <= "0000000000000000";
symbol_8(15) <= "0000000000000000";

symbol_9( 0) <= "0000000000000000";
symbol_9( 1) <= "0000000000000000";
symbol_9( 2) <= "0000000000000000";
symbol_9( 3) <= "0000111111110000";
symbol_9( 4) <= "0001111111111000";
symbol_9( 5) <= "0001100000011000";
symbol_9( 6) <= "0001100000011000";
symbol_9( 7) <= "0001111111111000";
symbol_9( 8) <= "0000111111111000";
symbol_9( 9) <= "0000000000011000";
symbol_9(10) <= "0001100000011000";
symbol_9(11) <= "0001111111111000";
symbol_9(12) <= "0000111111110000";
symbol_9(13) <= "0000000000000000";
symbol_9(14) <= "0000000000000000";
symbol_9(15) <= "0000000000000000";

begin
	dataOut <= symbol_player(to_integer(unsigned)address); --TODO
end Behavioral;
