library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use std.textio.ALL;
use IEEE.std_logic_textio.ALL;
use IEEE.Numeric_Std.All;

entity background is 
  Port ( clk       : in  std_logic;  -- 50 MHz clock
         reset     : in  std_logic;  -- reset signal
			background_rgb : in std_logic_vector(3 downto 0);
         AllX     : buffer std_logic_vector(639*479 downto 0);   -- horizontal coordinate
			AllXY    : buffer std_logic_vector(639*479 downto 0);
         AllY     : buffer std_logic_vector(479*638 downto 0) ); -- vertical coordinate
end background;

--add player position and check for collision. update maze based on collision

architecture Behavioral of background is
constant X_Center : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(320, 10);  --Center position on the X axis
constant Y_Center : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(240, 10);  --Center position on the Y axis
constant X_Min    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(0, 10);  --Leftmost point on the X axis
constant X_Max    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(639, 10);  --Rightmost point on the X axis
constant Y_Min    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(0, 10);   --Topmost point on the Y axis
constant Y_Max    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(479, 10);  --Bottommost point on the Y axis
signal X_border : std_logic_vector(639 downto 0);
signal Y_border : std_logic_vector(479 downto 0);

type array_molecule is array (29 downto 0) of std_logic_vector(159 downto 0); 
--type array_molecule is array (29 downto 0, 159 downto 0) of std_logic;
--add a new level flag to sensitivity list to check if new maze should be generated
signal maze_array : array_molecule :=
(
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111001100100010001000100010001000100010001000100010001000100010001000100010111111110010001000100010001000100010001000100010001000100010001000100010001000111111",
"1111001011111111111111111111111111110010111111111111111111111111111111110010111111110010111111111111111111111111111111110010111111111111111111111111111100101111",
"1111001011111111111111111111111111110010111111111111111111111111111111110010111111110010111111111111111111111111111111110010111111111111111111111111111100101111",
"1111001011111111111111111111111111110010111111111111111111111111111111110010111111110010111111111111111111111111111111110010111111111111111111111111111100101111",
"1111001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000101111",
"1111001011111111111111111111111111110010111111110010111111111111111111111111111111111111111111111111111111110010111111110010111111111111111111111111111100101111",
"1111001000100010001000100010001000100010111111110010111111111111111111111111111111111111111111111111111111110010111111110010001000100010001000100010001000101111",
"1111111111111111111111111111111111110010111111110010001000100010001000100010111111110010001000100010001000100010111111110010111111111111111111111111111111111111",
"1111111111111111111111111111111111110010111111111111111111111111111111110010111111110010111111111111111111111111111111110010111111111111111111111111111111111111",
"1111111111111111111111111111111111110010111111110010001000100010001000100010001000100010001000100010001000100010111111110010111111111111111111111111111111111111",
"1111111111111111111111111111111111110010111111110010111111111111111111111111000000001111111111111111111111110010111111110010111111111111111111111111111111111111",
"1111001000100010001000100010001000100010001000100010111100000000000000000000000000000000000000000000000011110010001000100010001000100010001000100010001000101111",
"1111111111111111111111111111111111110010111111110010111101000000000000000000000000000000000000000000010011110010111111110010111111111111111111111111111111111111",
"1111111111111111111111111111111111110010111111110010111111111111111111111111111111111111111111111111111111110010111111110010111111111111111111111111111111111111",
"1111111111111111111111111111111111110010111111110010001000100010001000100010001000100010001000100010001000100010111111110010111111111111111111111111111111111111",
"1111111111111111111111111111111111110010111111110010111111111111111111111111111111111111111111111111111111110010111111110010111111111111111111111111111111111111",
"1111001000100010001000100010001000100010001000100010001000100010001000100010111111110010001000100010001000100010001000100010001000100010001000100010001000101111",
"1111001011111111111111111111111111110010111111111111111111111111111111110010111111110010111111111111111111111111111111110010111111111111111111111111111100101111",
"1111001011111111111111111111111111110010111111111111111111111111111111110010111111110010111111111111111111111111111111110010111111111111111111111111111100101111",
"1111001000100010001000101111111111110010001000100010001000100010001000100010001000010010001000100010001000100010001000100010111111111111001000100010001000101111",
"1111111111111111111100101111111111110010111111110010111111111111111111111111111111111111111111111111111111110010111111110010111111111111001011111111111111111111",
"1111111111111111111100101111111111110010111111110010111111111111111111111111111111111111111111111111111111110010111111110010111111111111001011111111111111111111",
"1111001000100010001000100010001000100010111111110010001000100010001000100010111111110010001000100010001000100010111111110010001000100010001000100010001000101111",
"1111001011111111111111111111111111111111111111111111111111111111111111110010111111110010111111111111111111111111111111111111111111111111111111111111111100101111",
"1111001011111111111111111111111111111111111111111111111111111111111111110010111111110010111111111111111111111111111111111111111111111111111111111111111100101111",
"1111001100100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0001001000110100010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011110001001101010111100110111101111"
);

--begin
--TODO this code would potentially auto-generate a maze for each level
--background_rgb <= "000"; --TODO set to switches

--set_screen_borders: process(AllX, AllY)
--	variable I :
--			integer range 0 to 639;
--begin
--	set_Xborders: while (I<=639) loop
--		X_border(I) <= '1';
--		I := I + 1;
--	end loop set_Xborders;
--	
--	set_Yborders: while (I<=479) loop
--		Y_border(I) <= '1';
--		I := I + 1;
--	end loop set_Yborders;
--	
--	AllX(639 downto 0)<=X_border;
--	AllX(639*479 downto 639*478)<=X_border;
--	AllY(479 downto 0)<=Y_border;
--	AllY(479*639 downto 479*638)<=Y_border;
--	AllXY(639*479 downto 0)<=AllX(639*479 downto 0) OR AllY(639*479 downto 0);
----	report "Screen =" & integer'image(to_integer(TO_UNSIGNED((AllXY))));
----	write(AllXY(639*479 downto 0),"this should print the vector to screen");
--end process;

--print_to_screen: process (array_molecule)
--begin

--data <= ROM(to_integer(unsigned(addr)));
 
--end process;
end Behavioral;

--rectangle_on <= '1' when pixel_x >= 150 and pixel_x <= 250 and 
--                         pixel_y >= 100 and pixel_y <= 150 
--                  else '0';
--rectangle_rgb <= "111";9
--
--square_on <= '1' when pixel_x >= 350 and pixel_x <400 and 
--                      pixel_y >= 200 and pixel_y <250 
--              else '0';
--square_rgb <= "010";
--
---- Default value when no object is being displayed
--background_rgb <= "000";
--rgb_out <= rectangle_rgb when rectangle_on = '1' else
--             square_rgb when square_on = '1' else
--             background_rgb;